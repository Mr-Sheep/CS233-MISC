
module chopUpDigits_control (done, get_new, load_index, load_number, select_base, write, base, number_is_0, go, clk, reset);
	output done, get_new, load_index, load_number, select_base, write;
	input base, number_is_0, go;
	input clk, reset;

endmodule
